-- Copyright (C) 2017  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 17.1.0 Build 590 10/25/2017 SJ Lite Edition
-- Created on Mon May 13 14:08:48 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY DrinksFSM IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        V : IN STD_LOGIC := '0';
        C : IN STD_LOGIC := '0';
        drink : OUT STD_LOGIC
    );
END DrinksFSM;

ARCHITECTURE BEHAVIOR OF DrinksFSM IS
    TYPE type_fstate IS (E0,E1,E2,E3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,V,C)
    BEGIN
        IF (reset='0') THEN
            reg_fstate <= E0;
            drink <= '0';
        ELSE
            drink <= '0';
            CASE fstate IS
                WHEN E0 =>
                    IF ((NOT((C = '1')) AND NOT((V = '1')))) THEN
                        reg_fstate <= E0;
                    ELSIF ((NOT((C = '1')) AND (V = '1'))) THEN
                        reg_fstate <= E1;
                    ELSIF ((NOT((V = '1')) AND (C = '1'))) THEN
                        reg_fstate <= E2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E0;
                    END IF;

                    drink <= '0';
                WHEN E1 =>
                    IF ((NOT((C = '1')) AND NOT((V = '1')))) THEN
                        reg_fstate <= E1;
                    ELSIF ((NOT((C = '1')) AND (V = '1'))) THEN
                        reg_fstate <= E2;
                    ELSIF ((NOT((V = '1')) AND (C = '1'))) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E1;
                    END IF;

                    drink <= '0';
                WHEN E2 =>
                    IF ((NOT((C = '1')) AND NOT((V = '1')))) THEN
                        reg_fstate <= E2;
                    ELSIF (((C = '1') OR (V = '1'))) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E2;
                    END IF;

                    drink <= '0';
                WHEN E3 =>
                    reg_fstate <= E0;

                    drink <= '1';
                WHEN OTHERS => 
                    drink <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
